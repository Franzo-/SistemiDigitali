-- TOP LEVEL